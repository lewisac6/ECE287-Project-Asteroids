module title_spock_ascii #(
    parameter WIDTH  = 120,   
    parameter HEIGHT = 70,    
    parameter SCALE  = 8      
)(
    input  wire [9:0] pixel_x,
    input  wire [9:0] pixel_y,

    input  wire [9:0] origin_x,  
    input  wire [9:0] origin_y,

    output reg ascii_r,
    output reg ascii_g,
    output reg ascii_b
);

    reg [8*WIDTH-1:0] ascii [0:HEIGHT-1];
    integer i;

    initial begin
        ascii[0]  = "                     ..........................           ";
        ascii[1]  = "                 ...................................       ";
        ascii[2]  = "              .........................................    ";
        ascii[3]  = "            .............................................  ";
        ascii[4]  = "           ................................................ ";
        ascii[5]  = "          ..................................................";
        ascii[6]  = "         ....................................................";
        ascii[7]  = "         ......;%;%%%%%%%%%%%%%%%%%%%%%%%%%%%;%%..............";
        ascii[8]  = "         .....;%%%;;;;%%%%%%%%%%%%%%%%%%;;;;%%%%..............%";
        ascii[9]  = "         .....%%%%%%%%;;;%%%%%%%%%%%%;;;%%%%%%%%%............%%%";
        ascii[10] = "         /....%%%%%%%%%%%%;%%%%%%%%;%%%%%%%%%%%%%%..........;%%%";
        ascii[11] = "         //...%%%a@@`  '@%%//%%%%%%%%@`  '@@a%%%%%%........;%/%%";
        ascii[12] = "         //...%@@@@@aaa@@@%//%%%%%%@@@@aaa@@@@@%%%%%......%%/%%";
        ascii[13] = "         //...%%%%%%%%%%%%%//%%%%%%%%%%%%%%%%%%%%%%%%....%%/%%%";
        ascii[14] = "          //..%%%%%%%%%%%%//%%%%%%%%%%%%%%%%%%%%%%%%%...%%/%%%";
        ascii[15] = "           //.%%%%%%%%%%%%//%%%%%%%%%%%%%%%%%%%%%%%%%..%%/%%% ";
        ascii[16] = "            //%%%%%%%%%%%//%%%%%%%%%%%%%%%%%%%%%%%%%%..%/%%%  ";
        ascii[17] = "             ;%%%%%%%%%%%//%%%%%%%%%;/%%%%%%%%%%%%%%%.%%%     ";
        ascii[18] = "               %%%%%%%%%//%%%%%%%%%%%;/%%%%%%%%%%%%%%%%       ";
        ascii[19] = "                %%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%/        ";
        ascii[20] = "                 ;%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%//        ";
        ascii[21] = "                   %%%%%<<<<<<<<<<<<<<<<<%%%%%%%%%%;//        ";
        ascii[22] = "                    %%%%%<<<<<<<<<<<<<<<%%%%%%%%%%;///        ";
        ascii[23] = "                     %%%%%%%%%%%%%%%%%%%%%%%%%%%;/////        ";
        ascii[24] = "                      %%%%%%%%%%%%%%%%%%%%%%%%;///////.       ";
        ascii[25] = "                      /;%%%%%%%%%%%%%%%%%%%;////////....      ";
        ascii[26] = "                      ///;%%%%%%%%%%%%%%;////////.........    ";
        ascii[27] = "                    ...///////////////////////..............  ";
        ascii[28] = "                  ........////////////////................,;;,";
        ascii[29] = "               ,;............/////////.................,;;;;;;;;,";
        ascii[30] = "           ,;;;;;;,................................,;;;;;;;;;;;;;;,";
        ascii[31] = "       ,;;;;;;;;;;;;;,........................,;;;;;;;;;;;;;;;;;;;;";
        ascii[32] = "   ,;;;;;;;;;;;;;;;;;;;;;,................,;;;;;;;;;;;;;;;;;;;;;;;;";
        ascii[33] = " ,;;;;;;;;;;;;;;;;;;;;;;;;;;,.........,;;;;;;;;;;;;;;;;;;;;;;;;;;;; ";
        ascii[34] = ";;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;/#\\;;;;;;;;;;; ";
        ascii[35] = ";;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;/####\\;;;;;;;;; ";
        ascii[36] = ";;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;/#######\\;;;;;;; ";

        for (i = 37; i < HEIGHT; i = i + 1)
            ascii[i] = {8*WIDTH{1'b0}};
    end


    localparam integer CELL_W = SCALE;
    localparam integer CELL_H = SCALE;

    wire inside =
        (pixel_x >= origin_x) &&
        (pixel_x <  origin_x + WIDTH  * CELL_W) &&
        (pixel_y >= origin_y) &&
        (pixel_y <  origin_y + HEIGHT * CELL_H);

    wire [9:0] local_x = pixel_x - origin_x;
    wire [9:0] local_y = pixel_y - origin_y;

    // SCALE = 4 -> divide by 4 using >> 2
    wire [9:0] sx = local_x >> 2;  
    wire [9:0] sy = local_y >> 2; 

    reg [7:0] ch;

    always @* begin
        ascii_r = 1'b0;
        ascii_g = 1'b0;
        ascii_b = 1'b0;

        if (inside) begin
            ch = ascii[sy][(WIDTH-1-sx)*8 +: 8];
            if (ch != " " && ch != 8'd0) begin
                ascii_r = 1'b1;
                ascii_g = 1'b1;
                ascii_b = 1'b1;   
            end
        end
    end

endmodule
